library IEEE;
use IEEE.STD_LOGIC_1164.all;

package types_package is

	type cell_select_array is array (0 to 7) of std_logic_vector(7 downto 0);

end types_package;

package body types_package is
 
end types_package;
